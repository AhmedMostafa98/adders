`timescale 1ns / 1ps

module Lookahead(
						input [15:0] operand1, operand2,
						output Cout,
						output [15:0] Result
						);
	
	wire Cin;
	wire [15:0] P, G , C;
	wire [135:0] e;
	
	generate
		genvar i;
		for (i = 0; i<16; i = i + 1)
		begin : PG
			PG pg (.a(operand1[i]), .b(operand2[i]), .p(P[i]), .g(G[i]));
		end
	endgenerate
	
	//Cin = 0
	buf (Cin, 0);
	
	//C0 = G0 + P0.Cin
	and (e[0], P[0], Cin);
	or  (C[0], G[0], e[0]);
	
	//C1 = G1 + G0.P1 + P1.P0.Cin
	and (e[1], P[1], P[0], Cin);
	and (e[2], G[0], P[1]);
	or  (C[1], G[1], e[1], e[2]);
	
	//C2 = G2 + G1.P2 + G0.P2.P1 + P2.P1.P0.Cin
	and (e[3], P[2], P[1], P[0], Cin);
	and (e[4], G[0], P[2], P[1]);
	and (e[5], G[1], P[2]);
	or  (C[2], G[2], e[3], e[4] , e[5]);
	
	//C3 = G3 + G2.P3 + G1.P3.P2 + G0.P3.P2.P1 + P3.P2.P1.P0.Cin
	and (e[6], P[3], P[2], P[1], P[0], Cin);
	and (e[7], G[0], P[3], P[2], P[1]);
	and (e[8], G[1], P[3], P[2]);
	and (e[9], G[2], P[3]);
	or  (C[3], G[3], e[6], e[7], e[8] , e[9]);
	
	//C4 = G4 + G3.P4 + G2.P4.P3 + G1.P4.P3.P2 + G0.P4.P3.P2.P1 + P4.P3.P2.P1.P0.Cin
	and (e[10], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[11], G[0], P[4], P[3], P[2], P[1]);
	and (e[12], G[1], P[4], P[3], P[2]);
	and (e[13], G[2], P[4], P[3]);
	and (e[14], G[3], P[4]);
	or  (C[4], G[4], e[10], e[11], e[12] , e[13], e[14]);
	
	//C5 = G5 + G4.P5 + G3.P5.P4 + G2.P5.P4.P3 + G1.P5.P4.P3.P2 + G0.P5.P4.P3.P2.P1 + P5.P4.P3.P2.P1.P0.Cin
	and (e[15], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[16], G[0], P[5], P[4], P[3], P[2], P[1]);
	and (e[17], G[1], P[5], P[4], P[3], P[2]);
	and (e[18], G[2], P[5], P[4], P[3]);
	and (e[19], G[3], P[5], P[4]);
	and (e[20], G[4], P[5]);
	or  (C[5], G[5], e[15], e[16], e[17] , e[18], e[19], e[20]);
	
	//C6 = G6 + G5.P6 + G4.P6.P5 + G3.P6.P5.P4 + G2.P6.P5.P4.P3 + G1.P6.P5.P4.P3.P2 + G0.P6.P5.P4.P3.P2.P1 + P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[21], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[22], G[0], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[23], G[1], P[6], P[5], P[4], P[3], P[2]);
	and (e[24], G[2], P[6], P[5], P[4], P[3]);
	and (e[25], G[3], P[6], P[5], P[4]);
	and (e[26], G[4], P[6], P[5]);
	and (e[27], G[5], P[6]);
	or  (C[6], G[6], e[21], e[22], e[23] , e[24], e[25], e[26], e[27]);
	
	//C7 = G7 + G6.P7 + G5.P7.P6 + G4.P7.P6.P5 + G3.P7.P6.P5.P4 + G2.P7.P6.P5.P4.P3 + G1.P7.P6.P5.P4.P3.P2 + 
	//G0.P7.P6.P5.P4.P3.P2.P1 + P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[28], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[29], G[0], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[30], G[1], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[31], G[2], P[7], P[6], P[5], P[4], P[3]);
	and (e[32], G[3], P[7], P[6], P[5], P[4]);
	and (e[33], G[4], P[7], P[6], P[5]);
	and (e[34], G[5], P[7], P[6]);
	and (e[35], G[6], P[7]);
	or  (C[7], G[7], e[28], e[29], e[30] , e[31], e[32], e[33], e[34], e[35]);
	
	//C8 = G8 + G7.P8 + G6.P8.P7 + G5.P8.P7.P6 + G4.P8.P7.P6.P5 + G3.P8.P7.P6.P5.P4 + G2.P8.P7.P6.P5.P4.P3 + G1.P8.P7.P6.P5.P4.P3.P2 + 
	//G0.P8.P7.P6.P5.P4.P3.P2.P1 + P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[36], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[37], G[0], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[38], G[1], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[39], G[2], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[40], G[3], P[8], P[7], P[6], P[5], P[4]);
	and (e[41], G[4], P[8], P[7], P[6], P[5]);
	and (e[42], G[5], P[8], P[7], P[6]);
	and (e[43], G[6], P[8], P[7]);
	and (e[44], G[7], P[8]);
	or  (C[8], G[8], e[36], e[37], e[38] , e[39], e[40], e[41], e[42], e[43], e[44]);
	
	//C9 = G9 + G8.P9 + G7.P9.P8 + G6.P9.P8.P7 + G5.P9.P8.P7.P6 + G4.P9.P8.P7.P6.P5 + G3.P9.P8.P7.P6.P5.P4 + G2.P9.P8.P7.P6.P5.P4.P3 +
	//G1.P9.P8.P7.P6.P5.P4.P3.P2 + G0.P9.P8.P7.P6.P5.P4.P3.P2.P1 + P9.P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[45], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[46], G[0], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[47], G[1], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[48], G[2], P[9], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[49], G[3], P[9], P[8], P[7], P[6], P[5], P[4]);
	and (e[50], G[4], P[9], P[8], P[7], P[6], P[5]);
	and (e[51], G[5], P[9], P[8], P[7], P[6]);
	and (e[52], G[6], P[9], P[8], P[7]);
	and (e[53], G[7], P[9], P[8]);
	and (e[54], G[8], P[9]);
	or  (C[9], G[9], e[45], e[46], e[47] , e[48], e[49], e[50], e[51], e[52], e[53], e[54]);
	
	//C10 = G10 + G9.P10 + G8.P10.P9 + G7.P10.P9.P8 + G6.P10.P9.P8.P7 + G5.P10.P9.P8.P7.P6 + G4.P10.P9.P8.P7.P6.P5 +
	//G3.P10.P9.P8.P7.P6.P5.P4 + G2.P10.P9.P8.P7.P6.P5.P4.P3 + G1.P10.P9.P8.P7.P6.P5.P4.P3.P2 +
	//G0.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1 + P10.P9.P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[55], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[56], G[0], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[57], G[1], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[58], G[2], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[59], G[3], P[10], P[9], P[8], P[7], P[6], P[5], P[4]);
	and (e[60], G[4], P[10], P[9], P[8], P[7], P[6], P[5]);
	and (e[61], G[5], P[10], P[9], P[8], P[7], P[6]);
	and (e[62], G[6], P[10], P[9], P[8], P[7]);
	and (e[63], G[7], P[10], P[9], P[8]);
	and (e[64], G[8], P[10], P[9]);
	and (e[65], G[9], P[10]);
	or  (C[10], G[10], e[55], e[56], e[57] , e[58], e[59], e[60], e[61], e[62], e[63], e[64], e[65]);
	
	//C11 = G11 + G10.P11 + G9.P11.P10 + G8.P11.P10.P9 + G7.P11.P10.P9.P8 + G6.P11.P10.P9.P8.P7 + G5.P11.P10.P9.P8.P7.P6 + 
	//G4.P11.P10.P9.P8.P7.P6.P5 + G3.P11.P10.P9.P8.P7.P6.P5.P4 + G2.P11.P10.P9.P8.P7.P6.P5.P4.P3 + G1.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2 +
	//G0.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1 + P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[66], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[67], G[0], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[68], G[1], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[69], G[2], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[70], G[3], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4]);
	and (e[71], G[4], P[11], P[10], P[9], P[8], P[7], P[6], P[5]);
	and (e[72], G[5], P[11], P[10], P[9], P[8], P[7], P[6]);
	and (e[73], G[6], P[11], P[10], P[9], P[8], P[7]);
	and (e[74], G[7], P[11], P[10], P[9], P[8]);
	and (e[75], G[8], P[11], P[10], P[9]);
	and (e[76], G[9], P[11], P[10]);
	and (e[77], G[10], P[11]);
	or  (C[11], G[11], e[66], e[67], e[68] , e[69], e[70], e[71], e[72], e[73], e[74], e[75], e[76], e[77]);
	
	//C12 = G12 + G11.P12 + G10.P12.P11 + G9.P12.P11.P10 + G8.P12.P11.P10.P9 + G7.P12.P11.P10.P9.P8 + G6.P12.P11.P10.P9.P8.P7 + 
	//G5.P12.P11.P10.P9.P8.P7.P6 + G4.P12.P11.P10.P9.P8.P7.P6.P5 + G3.P12.P11.P10.P9.P8.P7.P6.P5.P4 +
	//G2.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3 + G1.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2 + G0.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1 + 
	//P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[78], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[79], G[0], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[80], G[1], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[81], G[2], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[82], G[3], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4]);
	and (e[83], G[4], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5]);
	and (e[84], G[5], P[12], P[11], P[10], P[9], P[8], P[7], P[6]);
	and (e[85], G[6], P[12], P[11], P[10], P[9], P[8], P[7]);
	and (e[86], G[7], P[12], P[11], P[10], P[9], P[8]);
	and (e[87], G[8], P[12], P[11], P[10], P[9]);
	and (e[88], G[9], P[12], P[11], P[10]);
	and (e[89], G[10], P[12], P[11]);
	and (e[90], G[11], P[12]);
	or  (C[12], G[12], e[78], e[79], e[80] , e[81], e[82], e[83], e[84], e[85], e[86], e[87], e[88], e[89], e[90]);
	
	//C13 = G13 + G12.P13 + G11.P13.P12 + G10.P13.P12.P11 + G9.P13.P12.P11.P10 + G8.P13.P12.P11.P10.P9 + G7.P13.P12.P11.P10.P9.P8 + 
	//G6.P13.P12.P11.P10.P9.P8.P7 + G5.P13.P12.P11.P10.P9.P8.P7.P6 + G4.P13.P12.P11.P10.P9.P8.P7.P6.P5 + 
	//G3.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4 + G2.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3 + G1.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2 + 
	//G0.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1 + P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[91], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[92], G[0], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[93], G[1], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[94], G[2], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[95], G[3], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4]);
	and (e[96], G[4], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5]);
	and (e[97], G[5], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6]);
	and (e[98], G[6], P[13], P[12], P[11], P[10], P[9], P[8], P[7]);
	and (e[99], G[7], P[13], P[12], P[11], P[10], P[9], P[8]);
	and (e[100], G[8], P[13], P[12], P[11], P[10], P[9]);
	and (e[101], G[9], P[13], P[12], P[11], P[10]);
	and (e[102], G[10], P[13], P[12], P[11]);
	and (e[103], G[11], P[13], P[12]);
	and (e[104], G[12], P[13]);
	or  (C[13], G[13], e[91], e[92], e[93] , e[94], e[95], e[96], e[97], e[98], e[99], e[100], e[101], e[102], e[103], e[104]);
	
	//C14 = G14 + G13.P14 + G12.P14.P13 + G11.P14.P13.P12 + G10.P14.P13.P12.P11 + G9.P14.P13.P12.P11.P10 + G8.P14.P13.P12.P11.P10.P9 + 
	//G7.P14.P13.P12.P11.P10.P9.P8 + G6.P14.P13.P12.P11.P10.P9.P8.P7 + G5.P14.P13.P12.P11.P10.P9.P8.P7.P6 + 
	//G4.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5 + G3.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4 + G2.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3 + 
	//G1.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2 + G0.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1 + 
	//P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[105], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[106], G[0], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[107], G[1], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[108], G[2], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[109], G[3], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4]);
	and (e[110], G[4], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5]);
	and (e[111], G[5], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6]);
	and (e[112], G[6], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7]);
	and (e[113], G[7], P[14], P[13], P[12], P[11], P[10], P[9], P[8]);
	and (e[114], G[8], P[14], P[13], P[12], P[11], P[10], P[9]);
	and (e[115], G[9], P[14], P[13], P[12], P[11], P[10]);
	and (e[116], G[10], P[14], P[13], P[12], P[11]);
	and (e[117], G[11], P[14], P[13], P[12]);
	and (e[118], G[12], P[14], P[13]);
	and (e[119], G[13], P[14]);
	or  (C[14], G[14], e[105], e[106], e[107] , e[108], e[109], e[110], e[111], e[112], e[113], e[114], e[115], e[116], e[117],
							 e[118], e[119]);
	
	//C15 = G15 + G14.P15 + G13.P15.P14 + G12.P15.P14.P13 + G11.P15.P14.P13.P12 + G10.P15.P14.P13.P12.P11 + G9.P15.P14.P13.P12.P11.P10 + 
	//G8.P15.P14.P13.P12.P11.P10.P9 + G7.P15.P14.P13.P12.P11.P10.P9.P8 + G6.P15.P14.P13.P12.P11.P10.P9.P8.P7 + 
	//G5.P15.P14.P13.P12.P11.P10.P9.P8.P7.P6 + G4.P15.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5 + G3.P15.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4 + 
	//G2.P15.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3 + G1.P15.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2 + 
	//G0.P15.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1 + P15.P14.P13.P12.P11.P10.P9.P8.P7.P6.P5.P4.P3.P2.P1.P0.Cin
	and (e[120], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1], P[0], Cin);
	and (e[121], G[0], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2], P[1]);
	and (e[122], G[1], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3], P[2]);
	and (e[123], G[2], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4], P[3]);
	and (e[124], G[3], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5], P[4]);
	and (e[125], G[4], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6], P[5]);
	and (e[126], G[5], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7], P[6]);
	and (e[127], G[6], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8], P[7]);
	and (e[128], G[7], P[15], P[14], P[13], P[12], P[11], P[10], P[9], P[8]);
	and (e[129], G[8], P[15], P[14], P[13], P[12], P[11], P[10], P[9]);
	and (e[130], G[9], P[15], P[14], P[13], P[12], P[11], P[10]);
	and (e[131], G[10], P[15], P[14], P[13], P[12], P[11]);
	and (e[132], G[11], P[15], P[14], P[13], P[12]);
	and (e[133], G[12], P[15], P[14], P[13]);
	and (e[134], G[13], P[15], P[14]);
	and (e[135], G[14], P[15]);
	or  (C[15], G[15], e[120], e[121], e[122] , e[123], e[124], e[125], e[126], e[127], e[128], e[129], e[130], e[131], e[132],
							 e[133], e[134], e[135]);
	
	
	//calculating sums
	xor (Result[0], P[0], Cin); // result = (A ^ B) . C;
	xor x[15:1] (Result [15:1], P[15:1], C[14:0]);
	buf (Cout, C[15]); // Cout = C15
	
endmodule
